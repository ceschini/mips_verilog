module logic_not(input A, output Y);
  assign Y = ~A;
endmodule