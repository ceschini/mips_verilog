module logic_and(input A, B, output Y);
  assign Y = A & B;
endmodule