module comparator (
  input [7:0] A,
   B,
   output [7:0] Amenor
);

  assign Amenor = ((~A[7] & B[7]) | (~(A[7] ^ B[7]) & (~A[6] & B[6]))
            | (~(A[7] ^ B[7]) & ~(A[6] ^ B[6]) & (~A[5] & B[5]))
            | (~(A[7] ^ B[7]) & ~(A[6] ^ B[6]) & ~(A[5] ^ B[5])
            & (~A[4] & B[4]))
            | (~(A[7] ^ B[7]) & ~(A[6] ^ B[6]) 
            & ~(A[5] ^ B[5]) & ~(A[4] ^ B[4])
            & (~A[3] & B[3]))
            | (~(A[7] ^ B[7]) & ~(A[6] ^ B[6]) 
            & ~(A[5] ^ B[5]) & ~(A[4] ^ B[4])
            & ~(A[3] ^ B[3])
            & (~A[2] & B[2]))
            | (~(A[7] ^ B[7]) & ~(A[6] ^ B[6]) 
            & ~(A[5] ^ B[5]) & ~(A[4] ^ B[4])
            & ~(A[3] ^ B[3]) & ~(A[2] ^ B[2])
            & (~A[1] & B[1]))
            | (~(A[7] ^ B[7]) & ~(A[6] ^ B[6]) 
            & ~(A[5] ^ B[5]) & ~(A[4] ^ B[4])
            & ~(A[3] ^ B[3]) & ~(A[2] ^ B[2])
            & ~(A[1] ^ B[1])
            & (~A[0] & B[0]))
                  ) ? 8'b11111111 : 8'b00000000;

endmodule
