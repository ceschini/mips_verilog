module logic_or(input A, B, output Y);
  assign Y = A | B;
endmodule